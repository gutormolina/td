LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_unsigned.all;

ENTITY counter IS
	PORT (
		load : IN std_logic;
		clk : IN std_logic;
		partidaS : IN std_logic_vector(5 downto 0);
		partidaM : IN std_logic_vector(5 downto 0);
		clear : IN std_logic;
		sentido : IN std_logic;
		hold : IN std_logic;
		fsel : IN std_logic;
		coutS : OUT std_logic_vector(13 downto 0);
		coutM : OUT std_logic_vector(13 downto 0)
	);
END counter;
ARCHITECTURE arch_counter OF counter IS
SIGNAL clkdiv : std_logic;
SIGNAL sigCountS, sigCountM: std_logic_vector(5 downto 0);
COMPONENT frequencyDivider
 PORT(
		clk50: IN std_logic;
		sel: IN std_logic;
		clk1: OUT std_logic
	);
END COMPONENT;
BEGIN
	fDiv: frequencyDivider
	PORT MAP(clk50 => clk, sel => fsel, clk1 => clkdiv);
	PROCESS(clear, clkdiv)
	VARIABLE countS, countM: std_logic_vector(5 downto 0);
		BEGIN
		IF clkdiv'EVENT AND clkdiv = '1' THEN
			IF clear = '1' THEN
				countS := "000000";
				countM := "000000";
			ELSIF load = '1' THEN
				countS := partidaS;
				countM := partidaM;
			ELSIF hold = '1' THEN
				countS := countS;
			ELSIF sentido = '1' THEN
				countS := countS - 1;
				IF countS = "000000" THEN
					countM := countM - 1;
					countS := "111011";
				END IF;
			ELSE
			   countS := countS + 1;
			END IF;
			IF countS = "111100" THEN
				countS := "000000";
				countM := countM + 1;
				end if;
		END IF;
		sigCountS <= countS;
		sigCountM <= countM;
	END PROCESS;
	
	WITH sigCountS SELECT
		coutS <=
			"00000010000001" WHEN "000000",
			"00000011001111" WHEN "000001",
			"00000010010010" WHEN "000010",
			"00000010000110" WHEN "000011",
			"00000011001100" WHEN "000100",
			"00000010100100" WHEN "000101",
			"00000010100000" WHEN "000110",
			"00000010001111" WHEN "000111",
			"00000010000000" WHEN "001000",
			"00000010000100" WHEN "001001",
			"10011110000001" WHEN "001010",
			"10011111001111" WHEN "001011",
			"10011110010010" WHEN "001100",
			"10011110000110" WHEN "001101",
			"10011111001100" WHEN "001110",
			"10011110100100" WHEN "001111",
			"10011110100000" WHEN "010000",
			"10011110001111" WHEN "010001",
			"10011110000000" WHEN "010010",
			"10011110000100" WHEN "010011",
			"00100100000001" WHEN "010100",
			"00100101001111" WHEN "010101",
			"00100100010010" WHEN "010110",
			"00100100000110" WHEN "010111",
			"00100101001100" WHEN "011000",
			"00100100100100" WHEN "011001",
			"00100100100000" WHEN "011010",
			"00100100001111" WHEN "011011",
			"00100100000000" WHEN "011100",
			"00100100000100" WHEN "011101",
			"00001100000001" WHEN "011110",
			"00001101001111" WHEN "011111",
			"00001100010010" WHEN "100000",
			"00001100000110" WHEN "100001",
			"00001101001100" WHEN "100010",
			"00001100100100" WHEN "100011",
			"00001100100000" WHEN "100100",
			"00001100001111" WHEN "100101",
			"00001100000000" WHEN "100110",
			"00001100000100" WHEN "100111",
			"10011000000001" WHEN "101000",
			"10011001001111" WHEN "101001",
			"10011000010010" WHEN "101010",
			"10011000000110" WHEN "101011",
			"10011001001100" WHEN "101100",
			"10011000100100" WHEN "101101",
			"10011000100000" WHEN "101110",
			"10011000001111" WHEN "101111",
			"10011000000000" WHEN "110000",
			"10011000000100" WHEN "110001",
			"01001000000001" WHEN "110010",
			"01001001001111" WHEN "110011",
			"01001000010010" WHEN "110100",
			"01001000000110" WHEN "110101",
			"01001001001100" WHEN "110110",
			"01001000100100" WHEN "110111",
			"01001000100000" WHEN "111000",
			"01001000001111" WHEN "111001",
			"01001000000000" WHEN "111010",
			"01001000000100" WHEN "111011",
			"11111101111110" WHEN OTHERS;
			
	WITH sigCountM SELECT
		coutM <=
			"00000010000001" WHEN "000000",
			"00000011001111" WHEN "000001",
			"00000010010010" WHEN "000010",
			"00000010000110" WHEN "000011",
			"00000011001100" WHEN "000100",
			"00000010100100" WHEN "000101",
			"00000010100000" WHEN "000110",
			"00000010001111" WHEN "000111",
			"00000010000000" WHEN "001000",
			"00000010000100" WHEN "001001",
			"10011110000001" WHEN "001010",
			"10011111001111" WHEN "001011",
			"10011110010010" WHEN "001100",
			"10011110000110" WHEN "001101",
			"10011111001100" WHEN "001110",
			"10011110100100" WHEN "001111",
			"10011110100000" WHEN "010000",
			"10011110001111" WHEN "010001",
			"10011110000000" WHEN "010010",
			"10011110000100" WHEN "010011",
			"00100100000001" WHEN "010100",
			"00100101001111" WHEN "010101",
			"00100100010010" WHEN "010110",
			"00100100000110" WHEN "010111",
			"00100101001100" WHEN "011000",
			"00100100100100" WHEN "011001",
			"00100100100000" WHEN "011010",
			"00100100001111" WHEN "011011",
			"00100100000000" WHEN "011100",
			"00100100000100" WHEN "011101",
			"00001100000001" WHEN "011110",
			"00001101001111" WHEN "011111",
			"00001100010010" WHEN "100000",
			"00001100000110" WHEN "100001",
			"00001101001100" WHEN "100010",
			"00001100100100" WHEN "100011",
			"00001100100000" WHEN "100100",
			"00001100001111" WHEN "100101",
			"00001100000000" WHEN "100110",
			"00001100000100" WHEN "100111",
			"10011000000001" WHEN "101000",
			"10011001001111" WHEN "101001",
			"10011000010010" WHEN "101010",
			"10011000000110" WHEN "101011",
			"10011001001100" WHEN "101100",
			"10011000100100" WHEN "101101",
			"10011000100000" WHEN "101110",
			"10011000001111" WHEN "101111",
			"10011000000000" WHEN "110000",
			"10011000000100" WHEN "110001",
			"01001000000001" WHEN "110010",
			"01001001001111" WHEN "110011",
			"01001000010010" WHEN "110100",
			"01001000000110" WHEN "110101",
			"01001001001100" WHEN "110110",
			"01001000100100" WHEN "110111",
			"01001000100000" WHEN "111000",
			"01001000001111" WHEN "111001",
			"01001000000000" WHEN "111010",
			"01001000000100" WHEN "111011",
			"11111101111110" WHEN OTHERS;
END arch_counter;